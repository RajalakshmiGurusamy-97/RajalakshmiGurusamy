//Public value only will get
class sample;
local int a;
protected int b;
int c;   //public
endclass
