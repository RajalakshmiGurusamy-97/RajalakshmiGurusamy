module tb;
parent p_inst;
   initial begin
   p_inst=new();
   p_inst.print();
   end
endmodule
